library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity transmitter is
    port (
        
    );
end entity transmitter;

architecture rtl of transmitter is
    
begin
    
    
    
end architecture rtl;